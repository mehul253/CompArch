
module test;
wire a;
assign a=1'b1;

reg b;
initial 
begin
    b=1'b1;
end
endmodule